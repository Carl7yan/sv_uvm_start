class test;
  env e0;

  function new();
    e0 = new;
  endfunction: new

  task run();
    e0.run;
  endtask: run
endclass: test
